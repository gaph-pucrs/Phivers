module Debug 
#(
    parameter PATH = "./"
)
(
    input  logic        clk_i,
    input  logic        rst_ni,

    input  logic        en_i,
    input  logic        we_i,
    input  logic [23:0] addr_i,
    input  logic [31:0] data_i
);

    /* @todo */

endmodule
